library ieee;
use ieee.std_logic_1164.all;

package lab_02_part_2_package is
   subtype part_2_vector is std_logic_vector;
end package lab_02_part_2_package;