library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package mas is
 type m is array(natural range<>) of integer;
end package mas;